`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//Testbench for top level
// 
//////////////////////////////////////////////////////////////////////////////////


module acsp_top_tb();


endmodule
